package typedefs;
    typedef 32 T; //number of timesteps cont.
    typedef 31 N_MAX; //number of max states w/o zero
    typedef 512 M_MAX; //number of max observations
    typedef 1024 INPUT_MAX;
endpackage